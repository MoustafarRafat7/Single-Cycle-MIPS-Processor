module Adder
(
input [31:0]input1,
input [31:0]input2,
output [31:0]out
);
assign out=input1+input2;
endmodule
